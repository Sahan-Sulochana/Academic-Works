

module test(

    );
endmodule
